module XOR (
    input wire A,
    input wire B,
    output wire F
);
    assign F = A ^ B;
endmodule