module NOT (
    input A,
    output F
);
    assign F = ~A;
endmodule